`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03.07.2023 22:18:56
// Design Name: 
// Module Name: LFadder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module LFadder(clk,A,B,cin,sum,cout);

//-------------------------------------PORTS DECLARATION----------------------------------//
input clk,cin;
input [15:0] A,B;
output reg [15:0] sum,cout;

//-------------------------------------INTERMEDIATE SIGNALS DECLARATION----------------------------------//
wire [15:0]G0,P0;
wire [7:0] G1,P1;
wire [6:0] G5,P5;
wire [3:0] G2,P2,G3,P3,G4,P4;
reg [15:0]G0_1,P0_1,G0_2,P0_2,G0_3,P0_3,G0_4,P0_4,G0_5,P0_5,P0_6;
reg [7:0] G1_2,P1_2,G1_3,P1_3,G1_4,P1_4,G1_5,P1_5;
reg [3:0] G2_3,P2_3,G2_4,P2_4,G2_5,P2_5,G3_4,P3_4,G3_5,P3_5,G4_5,P4_5;
reg [16:0]c1,c2,c3,c4,c5,c6;

//-------------------------------------FIRST STAGE G's AND P's GENERATION----------------------------------//

assign G0[0] = (A[0] & B[0]) | (cin & (A[0] | B[0])),
       G0[15:1] = A[15:1] & B[15:1];
     
assign P0 = A ^ B; 
       
//-------------------------------------FIRST STAGE G's AND P's REGISTERING----------------------------------//

always@(posedge clk)
    begin
        c1[0] <= cin;
        c1[1] <= G0[0];
        G0_1 <= G0;
        P0_1 <= P0;
    end 
    
//-------------------------------------SECOND STAGE G's AND P's GENERATION----------------------------------//
gp_gen i1_1(G0_1[1],G0_1[0],P0_1[1],P0_1[0],G1[0],P1[0]);
gp_gen i1_2(G0_1[3],G0_1[2],P0_1[3],P0_1[2],G1[1],P1[1]);
gp_gen i1_3(G0_1[5],G0_1[4],P0_1[5],P0_1[4],G1[2],P1[2]);
gp_gen i1_4(G0_1[7],G0_1[6],P0_1[7],P0_1[6],G1[3],P1[3]);
gp_gen i1_5(G0_1[9],G0_1[8],P0_1[9],P0_1[8],G1[4],P1[4]);
gp_gen i1_6(G0_1[11],G0_1[10],P0_1[11],P0_1[10],G1[5],P1[5]);
gp_gen i1_7(G0_1[13],G0_1[12],P0_1[13],P0_1[12],G1[6],P1[6]);
gp_gen i1_8(G0_1[15],G0_1[14],P0_1[15],P0_1[14],G1[7],P1[7]);

//-------------------------------------SECOND STAGE G's AND P's REGISTERING----------------------------------//

always@(posedge clk)
    begin
        c2[0] <= c1[0];
        c2[1] <= c1[1];
        c2[2] <= G1[0];
        G0_2 <= G0_1;
        P0_2 <= P0_1;
        G1_2 <= G1;
        P1_2 <= P1;
    end 
    
 //-------------------------------------THIRD STAGE G's AND P's GENERATION----------------------------------//   
 gp_gen i2_1(G1_2[1],G1_2[0],P1_2[1],P1_2[0],G2[0],P2[0]);
 gp_gen i2_2(G1_2[3],G1_2[2],P1_2[3],P1_2[2],G2[1],P2[1]);
 gp_gen i2_3(G1_2[5],G1_2[4],P1_2[5],P1_2[4],G2[2],P2[2]);
 gp_gen i2_4(G1_2[7],G1_2[6],P1_2[7],P1_2[6],G2[3],P2[3]);
 
 //-------------------------------------THIRD STAGE G's AND P's REGISTERING----------------------------------//

always@(posedge clk)
    begin
        c3[0] <= c2[0];
        c3[1] <= c2[1];
        c3[2] <= c2[2];
        c3[4] <= G2[0];
        G0_3 <= G0_2;
        P0_3 <= P0_2;
        G1_3 <= G1_2;
        P1_3 <= P1_2;
        G2_3 <= G2;
        P2_3 <= P2;
    end 
    
 //-------------------------------------FOURTH STAGE G's AND P's GENERATION----------------------------------//   
 gp_gen i3_1(G1_3[2],G2_3[0],P1_3[2],P2_3[0],G3[0],P3[0]);
 gp_gen i3_2(G2_3[1],G2_3[0],P2_3[1],P2_3[0],G3[1],P3[1]);
 gp_gen i3_3(G1_3[6],G2_3[2],P1_3[6],P2_3[2],G3[2],P3[2]);
 gp_gen i3_4(G2_3[3],G2_3[2],P2_3[3],P2_3[2],G3[3],P3[3]);
 
 //-------------------------------------FOURTH STAGE G's AND P's REGISTERING----------------------------------//

always@(posedge clk)
    begin
        c4[0] <= c3[0];
        c4[1] <= c3[1];
        c4[2] <= c3[2];
        c4[4] <= c3[4];
        c4[6] <= G3[0];
        c4[8] <= G3[1];
        G0_4 <= G0_3;
        P0_4 <= P0_3;
        G1_4 <= G1_3;
        P1_4 <= P1_3;
        G2_4 <= G2_3;
        P2_4 <= P2_3;
        G3_4 <= G3;
        P3_4 <= P3;
    end   
    
 //-------------------------------------FIFTH STAGE G's AND P's GENERATION----------------------------------//   
 gp_gen i4_1(G1_4[4],G3_4[1],P1_4[4],P3_4[1],G4[0],P4[0]);
 gp_gen i4_2(G2_4[2],G3_4[1],P2_4[2],P3_4[1],G4[1],P4[1]);
 gp_gen i4_3(G3_4[2],G3_4[1],P3_4[2],P3_4[1],G4[2],P4[2]);
 gp_gen i4_4(G3_4[3],G3_4[1],P3_4[3],P3_4[1],G4[3],P4[3]);
 
 //-------------------------------------FIFTH STAGE G's AND P's REGISTERING----------------------------------//

always@(posedge clk)
    begin
        c5[0] <= c4[0];
        c5[1] <= c4[1];
        c5[2] <= c4[2];
        c5[4] <= c4[4];
        c5[6] <= c4[6];
        c5[8] <= c4[8];
        c5[10] <= G4[0];
        c5[12] <= G4[1];
        c5[14] <= G4[2];
        c5[16] <= G4[3];
        G0_5 <= G0_4;
        P0_5 <= P0_4;
        G1_5 <= G1_4;
        P1_5 <= P1_4;
        G2_5 <= G2_4;
        P2_5 <= P2_4;
        G3_5 <= G3_4;
        P3_5 <= P3_4;
        G4_5 <= G4;
        P4_5 <= P4;
    end  
    
 //-------------------------------------SIXTH STAGE G's AND P's GENERATION----------------------------------//   
 gp_gen i5_1(G0_5[2],G1_5[0],P0_5[0],P1_5[0],G5[0],P5[0]);
 gp_gen i5_2(G0_5[4],G2_5[0],P0_5[4],P2_5[0],G5[1],P5[1]);
 gp_gen i5_3(G0_5[6],G3_5[0],P0_5[6],P3_5[0],G5[2],P5[2]);
 gp_gen i5_4(G0_5[8],G3_5[1],P0_5[8],P3_5[1],G5[3],P5[3]);
 gp_gen i5_5(G0_5[10],G4_5[0],P0_5[10],P4_5[0],G5[4],P5[4]);
 gp_gen i5_6(G0_5[12],G4_5[1],P0_5[12],P4_5[1],G5[5],P5[5]);
 gp_gen i5_7(G0_5[14],G4_5[2],P0_5[14],P4_5[2],G5[6],P5[6]);
 
 //-------------------------------------SIXTH STAGE G's AND P's REGISTERING----------------------------------//

always@(posedge clk)
    begin
        c6[0] <= c5[0];
        c6[1] <= c5[1];
        c6[2] <= c5[2];
        c6[4] <= c5[4];
        c6[6] <= c5[6];
        c6[8] <= c5[8];
        c6[10] <= c5[10];
        c6[12] <= c5[12];
        c6[14] <= c5[14];
        c6[16] <= c5[16];
        c6[3] <= G5[0];
        c6[5] <= G5[1];
        c6[7] <= G5[2];
        c6[9] <= G5[3];
        c6[11] <= G5[4];
        c6[13] <= G5[5];
        c6[15] <= G5[6];
        P0_6 <= P0_5;
    end  
    
//-------------------------------------SUM CALCULATION----------------------------------// 
always@(posedge clk)
    begin
        sum <= c6[15:0] ^ P0_6;
        cout <= c6[16];
    end             
endmodule