`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02.07.2023 11:09:49
// Design Name: 
// Module Name: BKadder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module BKadder(A,B,Cin,clk,Sum,Cout);
input [15:0] A,B;
input Cin,clk;
output reg [15:0] Sum;
output reg Cout;

wire [15:0] P0,G0;
wire [7:0] P1,G1;
wire [3:0] P2,G2;
wire [1:0] P3,G3;
wire P4,G4;
reg [15:0] P0_1,G0_1,P0_2,G0_2,P0_3,G0_3,P0_4,G0_4,P0_5,G0_5,P0_6,G0_6,P0_7;
reg [7:0] P1_2,G1_2,P1_3,G1_3,P1_4,G1_4,G1_5,P1_5;
reg [3:0] P2_3,G2_3,P2_4,G2_4;
reg [1:0] G3_4,P3_4;
reg [15:0] C1,C2,C3,C4,C5,C6,C7;
reg Cout5,Cout6,Cout7;


/* ============ 1st stage ============================== */

assign G0[0]= (A[0] & B[0]) | (Cin & (A[0] | B[0])),
	   G0[1]= A[1] & B[1],
	   G0[2]= A[2] & B[2],
	   G0[3]= A[3] & B[3],
	   G0[4]= A[4] & B[4],
	   G0[5]= A[5] & B[5],
	   G0[6]= A[6] & B[6],
	   G0[7]= A[7] & B[7],
	   G0[8]= A[8] & B[8],
	   G0[9]= A[9] & B[9],
	   G0[10]= A[10] & B[10],
	   G0[11]= A[11] & B[11],
	   G0[12]= A[12] & B[12],
	   G0[13]= A[13] & B[13],
	   G0[14]= A[14] & B[14],
	   G0[15]= A[15] & B[15];
					

assign P0[0]= A[0] ^ B[0],
	   P0[1]= A[1] ^ B[1],
	   P0[2]= A[2] ^ B[2],
	   P0[3]= A[3] ^ B[3],
	   P0[4]= A[4] ^ B[4],
	   P0[5]= A[5] ^ B[5],
	   P0[6]= A[6] ^ B[6],
	   P0[7]= A[7] ^ B[7],
	   P0[8]= A[8] ^ B[8],
	   P0[9]= A[9] ^ B[9],
	   P0[10]= A[10] ^ B[10],
	   P0[11]= A[11] ^ B[11],
	   P0[12]= A[12] ^ B[12],
	   P0[13]= A[13] ^ B[13],
	   P0[14]= A[14] ^ B[14],
	   P0[15]= A[15] ^ B[15];
always@(posedge clk)
begin
    C1[1] <= G0[0];
    C1[0] <= Cin;
    P0_1 <= P0;
    G0_1 <= G0;
end

//=========2nd set=====================// 
assign P1[0]=P0_1[1] & P0_1[0],
	   P1[1]=P0_1[3] & P0_1[2],
	   P1[2]=P0_1[5] & P0_1[4],
	   P1[3]=P0_1[7] & P0_1[6],
	   P1[4]=P0_1[9] & P0_1[8],
	   P1[5]=P0_1[11] & P0_1[10],
	   P1[6]=P0_1[13] & P0_1[12],
	   P1[7]=P0_1[15] & P0_1[14];

assign G1[0]=G0_1[1]|(P0_1[1] & G0_1[0]),
	   G1[1]=G0_1[3]|(P0_1[3] & G0_1[2]),
	   G1[2]=G0_1[5]|(P0_1[5] & G0_1[4]),
	   G1[3]=G0_1[7]|(P0_1[7] & G0_1[6]),
	   G1[4]=G0_1[9]|(P0_1[9] & G0_1[8]),
	   G1[5]=G0_1[11]|(P0_1[11] & G0_1[10]),
	   G1[6]=G0_1[13]|(P0_1[13] & G0_1[12]),
	   G1[7]=G0_1[15]|(P0_1[15] & G0_1[14]);

always@(posedge clk)
begin
C2[1] <= C1[1];
C2[2] <= G1[0];
C2[0] <= C1[0];
P0_2 <= P0_1;
G0_2 <= G0_1;
P1_2 <= P1;
G1_2 <= G1;
end

// ============= 3rd set ========================//
assign P2[0]=P1_2[1] & P1_2[0],
	   P2[1]=P1_2[3] & P1_2[2],
	   P2[2]=P1_2[5] & P1_2[4],
	   P2[3]=P1_2[7] & P1_2[6];



assign G2[0] =G1_2[1]| (P1_2[1] &  G1_2[0]),
	   G2[1] =G1_2[3]| (P1_2[3] &  G1_2[2]),
	   G2[2]=G1_2[5]|(P1_2[5] & G1_2[4]),
	   G2[3]=G1_2[7]|(P1_2[7] & G1_2[6]);
	   
	   
always@(posedge clk)
begin
C3[4] <= G2[0];
C3[3] <= G0_2[2] | (P0_2[2] & C2[2]);
C3[1] <= C2[1];
C3[2] <= C2[2];
C3[0] <= C2[0];
P0_3 <= P0_2;
G0_3 <= G0_2;
P1_3 <= P1_2;
G1_3 <= G1_2;
P2_3 <= P2;
G2_3 <= G2;
end

//=================4th stage set==========//

assign P3[0]=P2_3[1] & P2_3[0],
	   P3[1]=P2_3[3] & P2_3[2];

assign G3[0]=G2_3[1]|(P2_3[1] & G2_3[0]),
	   G3[1]=G2_3[3]|(P2_3[3] & G2_3[2]);

always@(posedge clk)
begin
C4[8] <= G3[0];
C4[5] <= G0_3[4]| (P0_3[4]&C3[4]);
C4[6] <= G1_3[2]| (P1_3[2]& C3[4]);

C4[4] <= C3[4];
C4[3] <= C3[3];
C4[2] <= C3[2];
C4[1] <= C3[1];
C4[0] <= C3[0];

P0_4 <= P0_3;
G0_4 <= G0_3;
P1_4 <= P1_3;
G1_4 <= G1_3;
P2_4 <= P2_3;
G2_4 <= G2_3;
G3_4 <= G3;
P3_4 <= P3;

end

// ==========5th stage ==============//

assign P4= P3_4[1] & P3_4[0];

assign G4 = G3_4[1]|(P3_4[1] & G3_4[0]);

always@(posedge clk)
begin 
Cout5 <= G4;
C5[7] <= G0_4[6]| (P0_4[6] & C4[6]);
C5[9] <= G0_4[8]| (P0_4[8] & C4[8]);
C5[10] <= G1_4[4]| (P1_4[4] & C4[8]);
C5[12] <= G2_4[2]| (P2_4[2] & C4[8]);

C5[8] <= C4[8];
C5[5] <= C4[5];
C5[6] <= C4[6];
C5[4] <= C4[4];
C5[3] <= C4[3];
C5[2] <= C4[2];
C5[1] <= C4[1];
C5[0] <= C4[0];

P0_5 <= P0_4;
G0_5 <= G0_4;
P1_5 <= P1_4;
G1_5 <= G1_4;
end

// =========== 6th stage ==============//
always@(posedge clk)
begin
C6[11] <= G0_5[10]| (P0_5[10]&C5[10]);
C6[13] <= G0_5[12]| (P0_5[12]&C5[12]);
C6[14] <= G1_5[6]| (P1_5[6]&C5[12]);


C6[12] <= C5[12];
C6[10] <= C5[10];
C6[9] <= C5[9];
C6[8] <= C5[8];
C6[7] <= C5[7];
C6[5] <= C5[5];
C6[6] <= C5[6];
C6[4] <= C5[4];
C6[3] <= C5[3];
C6[2] <= C5[2];
C6[1] <= C5[1];
C6[0] <= C5[0];
Cout6 <= Cout5;

P0_6 <= P0_5;
G0_6 <= G0_5;
end

//=========== 7th stage ============//
always@(posedge clk)
begin
C7[15] <= G0_6[14]| (P0_6[14]&C6[14]);
C7[14] <= C6[14];
C7[13] <= C6[13];
C7[12] <= C6[12];
C7[11] <= C6[11];
C7[10] <= C6[10];
C7[9] <= C6[9];
C7[8] <= C6[8];
C7[7] <= C6[7];
C7[6] <= C6[6];
C7[5] <= C6[5];
C7[4] <= C6[4];
C7[3] <= C6[3];
C7[2] <= C6[2];
C7[1] <= C6[1];
C7[0] <= C6[0];
Cout7 <= Cout6;

P0_7 <= P0_6;
end

//========= 8th stage ============//
always@(posedge clk)
begin
/*C8[15]=C7[15];
C8[14]=C7[14];
C8[13]=C7[13];
C8[12]=C7[12];
C8[11]=C7[11];
C8[10]=C7[10];
C8[9]=C6[9];
C8[8]=C7[8];
C8[7]=C7[7];
C8[6]=C7[6];
C8[5]=C7[5];
C8[4]=C7[4];
C8[3]=C7[3];
C8[2]=C7[2];
C8[1]=C7[1];
C8[0]=C7[0];
P0_8=P0_7;*/
Cout <= Cout7;

Sum[0] <= P0_7[0]^C7[0];
Sum[1] <= P0_7[1]^C7[1];
Sum[2] <= P0_7[2]^C7[2];
Sum[3] <= P0_7[3]^C7[3];
Sum[4] <= P0_7[4]^C7[4];
Sum[5] <= P0_7[5]^C7[5];
Sum[6] <= P0_7[6]^C7[6];
Sum[7] <= P0_7[7]^C7[7];
Sum[8] <= P0_7[8]^C7[8];
Sum[9] <= P0_7[9]^C7[9];
Sum[10] <= P0_7[10]^C7[10];
Sum[11] <= P0_7[11]^C7[11];
Sum[12] <= P0_7[12]^C7[12];
Sum[13] <= P0_7[13]^C7[13];
Sum[14] <= P0_7[14]^C7[14];
Sum[15] <= P0_7[14]^C7[15];
end

endmodule


