`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03.07.2023 23:29:54
// Design Name: 
// Module Name: HCadder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module HCadder(A,B,Cin,clk,Sum,Cout);
input [15:0] A,B;
input Cin,clk;
output reg [15:0] Sum;
output reg Cout;

reg  Cin_0,Cin_1,Cin_2,Cin_3,Cin_4,Cin_5;

wire [15:0] G0,P0;
reg [15:0] G0_0,G0_1,G0_2,G0_3,G0_4,P0_0,P0_1,P0_2,P0_3,P0_4,P0_5;
//================== 0 stage  =========//

assign G0[0]= (A[0] & B[0])| (Cin & (A[0] | B[0])),
       G0[15:1]=A[15:1] & B[15:1],
	   P0 = A ^ B;
	   
always@(posedge clk)
begin
G0_0 <= G0;
P0_0 <= P0;
Cin_0 <= Cin;
end 

//========================  1st stage ==========================//
wire [7:0] G1,P1;
reg [7:0] G1_1,P1_1;

assign G1[0]=G0_0[1] | (P0_0[1] & G0_0[0]),
       G1[1]=G0_0[3] | (P0_0[3] & G0_0[2]),
	   G1[2]=G0_0[5] | (P0_0[5] & G0_0[4]),
	   G1[3]=G0_0[7] | (P0_0[7] & G0_0[6]),
	   G1[4]=G0_0[9] | (P0_0[9] & G0_0[8]),
       G1[5]=G0_0[11] | (P0_0[11] & G0_0[10]),
	   G1[6]=G0_0[13] | (P0_0[13] & G0_0[12]),
	   G1[7]=G0_0[15] | (P0_0[15] & G0_0[14]);
	   
assign P1[0] = P0_0[1] & P0_0[0],
       P1[1] = P0_0[3] & P0_0[2],
	   P1[2] = P0_0[5] & P0_0[4],
       P1[3] = P0_0[7] & P0_0[6],
	   P1[4] = P0_0[9] & P0_0[8],
       P1[5] = P0_0[11] & P0_0[10],
	   P1[6] = P0_0[13] & P0_0[12],
       P1[7] = P0_0[15] & P0_0[14];
	   
always@(posedge clk)
begin

P1_1 <= P1;
G1_1 <= G1;

G0_1 <= G0_0 ;
P0_1 <= P0_0 ;
Cin_1 <= Cin_0;

end

//=====================  2nd stage  ==================//
wire [6:0] G2,P2;
reg [6:0] G2_2,P2_2;
reg G1_2,P1_2,G1_3,P1_3,G1_4,P1_4;

assign G2[6:0] = G1_1[7:1] | (P1_1[7:1] & G1_1[6:0]);
assign  P2[6:0] = P1_1[7:1] & P1_1[6:0];

always@(posedge clk)
begin
G2_2 <= G2;
P2_2 <= P2;

G1_2 <= G1_1[0];
P1_2 <= P1_1[0];

G0_2 <= G0_1;
P0_2 <= P0_1;
Cin_2 <= Cin_1;

end

//======================== 3rd stage ===================//
wire [5:0] G3,P3;
reg [5:0] G3_3,P3_3;
reg G2_3,P2_3,G2_4,P2_4;

assign G3[5:1] = G2_2[6:2] | (P2_2[6:2] & G2_2[4:0]),
       G3[0] = G2_2[1] | (P2_2[1] & G1_2);
	   
assign P3[5:1] = P2_2[6:2] & P2_2[4:0],
	   P3[0] = P2_2[1] & P1_2;
	   
always@(posedge clk)
begin
G3_3 <= G3;
P3_3 <= P3;

G2_3 <= G2_2[0];
P2_3 <= P2_2[0];

G1_3 <= G1_2;
P1_3 <= P1_2;

G0_3 <= G0_2;
P0_3 <= P0_2;
Cin_3 <= Cin_2;
end

//=========================  4th stage ==========================//
wire [3:0] P4,G4;
reg [3:0] P4_4,G4_4;
reg P3_4_0,P3_4_1,G3_4_0,G3_4_1;


assign G4[0]= G3_3[2] | (P3_3[2] & G1_3),
       G4[1]= G3_3[3] | (P3_3[3] & G2_3),
	   G4[2]= G3_3[4] | (P3_3[4] & G3_3[0]),
	   G4[3]= G3_3[5] | (P3_3[5] & G3_3[1]);
	   
assign P4[0]=P3_3[2] & P1_3,
       P4[1]=P3_3[3] & P2_3,
	   P4[2]=P3_3[4] & P3_3[0],
	   P4[3]=P3_3[5] & P3_3[1];
	   
always@(posedge clk)
begin
P4_4 <= P4;
G4_4 <= G4;

G3_4_0 <= G3_3[0];
G3_4_1 <= G3_3[1];
P3_4_0 <= P3_3[0];
P3_4_1 <= P3_3[1];

G2_4  <= G2_3;
P2_4  <= P2_3;
 
G1_4  <= G1_3;
P1_4  <= P1_3;
 
G0_4  <= G0_3;
P0_4  <= P0_3; 
Cin_4 <= Cin_3;

end


// =========================  5th stage =================================//

wire [6:0] G5;
reg [15:0] G5_5;

assign G5[0]= G0_4[2] | (P0_4[2] & G1_4),
       G5[1]= G0_4[4] | (P0_4[4] & G2_4),
	   G5[2]= G0_4[6] | (P0_4[6] & G3_4_0),
	   G5[3]= G0_4[8] | (P0_4[8] & G3_4_1),
	   G5[4]= G0_4[10] | (P0_4[10] & G4_4[0]),
       G5[5]= G0_4[12] | (P0_4[12] & G4_4[1]),
	   G5[6]= G0_4[14] | (P0_4[14] & G4_4[2]);
	   
always@(posedge clk)
begin
G5_5[0] <= G0_4[0];
G5_5[1] <= G1_4;
G5_5[2] <= G5[0];
G5_5[3] <= G2_4;
G5_5[4] <= G5[1];
G5_5[5] <= G3_4_0;
G5_5[6] <= G5[2];
G5_5[7] <= G3_4_1;
G5_5[8] <= G5[3];
G5_5[9] <= G4_4[0];
G5_5[10] <= G5[4];
G5_5[11] <= G4_4[1];
G5_5[12] <= G5[5];
G5_5[13] <= G4_4[2];
G5_5[14] <= G5[6];
G5_5[15] <= G4_4[3];

P0_5  <= P0_4; 
Cin_5 <= Cin_4;
end

// =============== 6th stage sum calculation =========//

always@(posedge clk)
begin
Cout <= G5_5[15];
Sum[0] <= P0_5[0] ^ Cin_5;
Sum[15:1] <= P0_5[15:1] ^ G5_5[14:0];
end

endmodule


	   
	   
